module aha(a,b,s);
input a,b;
output s; 

assign s = a ^ b;

endmodule
